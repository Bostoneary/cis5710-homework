/* INSERT NAME AND PENNKEY HERE */
// NAME:Zhiye Zhang
// PENNKEY:zhiyez

`timescale 1ns / 1ns

// quotient = dividend / divisor

module divider_unsigned (
    input  wire [31:0] i_dividend,
    input  wire [31:0] i_divisor,
    output wire [31:0] o_remainder,
    output wire [31:0] o_quotient
);

    // TODO: your code here

endmodule


module divu_1iter (
    input  wire [31:0] i_dividend,
    input  wire [31:0] i_divisor,
    input  wire [31:0] i_remainder,
    input  wire [31:0] i_quotient,
    output wire [31:0] o_dividend,
    output wire [31:0] o_remainder,
    output wire [31:0] o_quotient
);
  /*
    for (int i = 0; i < 32; i++) {
        remainder = (remainder << 1) | ((dividend >> 31) & 0x1);
        if (remainder < divisor) {
            quotient = (quotient << 1);
        } else {
            quotient = (quotient << 1) | 0x1;
            remainder = remainder - divisor;
        }
        dividend = dividend << 1;
    }
    */
    logic [31:0] remainder_cmp;

    // TODO: your code here
    assign remainder_cmp=(i_remainder<<1)|((i_dividend>>31)&32'b1);
    assign o_remainder=(remainder_cmp>=i_divisor)?(remainder_cmp-i_divisor):remainder_cmp;
    assign o_quotient=(remainder_cmp>=i_divisor)?((i_quotient<<1)&32'b1):(i_quotient<<1);
    assign o_dividend=i_dividend<<1;

endmodule
